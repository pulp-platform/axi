module axi_rt_unit #()();

endmodule
