// Copyright 2020 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Authors:
// - Matheus Cavalcante <matheusd@iis.ee.ethz.ch>

// NOTE: The upsizer does not support WRAP bursts, and will answer with SLVERR
// upon receiving a burst of such type. In addition to that, the downsizer also
// does not support FIXED bursts with incoming axlen != 0.

module axi_dw_converter #(
    parameter int unsigned MaxReads         = 1    , // Number of outstanding reads
    parameter int unsigned SlvPortDataWidth = 8    , // Data width of the slv port
    parameter int unsigned MstPortDataWidth = 8    , // Data width of the mst port
    parameter int unsigned AddrWidth        = 1    , // Address width
    parameter int unsigned IdWidth          = 1    , // ID width
    parameter type aw_chan_t                = logic, // AW Channel Type
    parameter type mst_w_chan_t             = logic, //  W Channel Type for the mst port
    parameter type slv_w_chan_t             = logic, //  W Channel Type for the slv port
    parameter type b_chan_t                 = logic, //  B Channel Type
    parameter type ar_chan_t                = logic, // AR Channel Type
    parameter type mst_r_chan_t             = logic, //  R Channel Type for the mst port
    parameter type slv_r_chan_t             = logic, //  R Channel Type for the slv port
    parameter type mst_port_axi_req_t       = logic, // AXI Request Type for mst ports
    parameter type mst_port_axi_rsp_t       = logic, // AXI Response Type for mst ports
    parameter type slv_port_axi_req_t       = logic, // AXI Request Type for slv ports
    parameter type slv_port_axi_rsp_t       = logic  // AXI Response Type for slv ports
  ) (
    input  logic              clk_i,
    input  logic              rst_ni,
    // Slave interface
    input  slv_port_axi_req_t slv_req_i,
    output slv_port_axi_rsp_t slv_rsp_o,
    // Master interface
    output mst_port_axi_req_t mst_req_o,
    input  mst_port_axi_rsp_t mst_rsp_i
  );

  if (MstPortDataWidth == SlvPortDataWidth) begin: gen_no_dw_conversion
    assign mst_req_o = slv_req_i ;
    assign slv_rsp_o = mst_rsp_i;
  end : gen_no_dw_conversion

  if (MstPortDataWidth > SlvPortDataWidth) begin: gen_dw_upsize
    axi_dw_upsizer #(
      .MaxReads           (MaxReads        ),
      .SlvPortDataWidth   (SlvPortDataWidth),
      .MstPortDataWidth   (MstPortDataWidth),
      .AddrWidth          (AddrWidth       ),
      .IdWidth            (IdWidth         ),
      .aw_chan_t          (aw_chan_t          ),
      .mst_w_chan_t       (mst_w_chan_t       ),
      .slv_w_chan_t       (slv_w_chan_t       ),
      .b_chan_t           (b_chan_t           ),
      .ar_chan_t          (ar_chan_t          ),
      .mst_r_chan_t       (mst_r_chan_t       ),
      .slv_r_chan_t       (slv_r_chan_t       ),
      .mst_port_axi_req_t (mst_port_axi_req_t ),
      .mst_port_axi_rsp_t (mst_port_axi_rsp_t ),
      .slv_port_axi_req_t (slv_port_axi_req_t ),
      .slv_port_axi_rsp_t (slv_port_axi_rsp_t )
    ) i_axi_dw_upsizer (
      .clk_i     (clk_i    ),
      .rst_ni    (rst_ni   ),
      // Slave interface
      .slv_req_i (slv_req_i),
      .slv_rsp_o (slv_rsp_o),
      // Master interface
      .mst_req_o (mst_req_o),
      .mst_rsp_i (mst_rsp_i)
    );
  end : gen_dw_upsize

  if (MstPortDataWidth < SlvPortDataWidth) begin: gen_dw_downsize
    axi_dw_downsizer #(
      .MaxReads           (MaxReads        ),
      .SlvPortDataWidth   (SlvPortDataWidth),
      .MstPortDataWidth   (MstPortDataWidth),
      .AddrWidth          (AddrWidth       ),
      .IdWidth            (IdWidth         ),
      .aw_chan_t          (aw_chan_t          ),
      .mst_w_chan_t       (mst_w_chan_t       ),
      .slv_w_chan_t       (slv_w_chan_t       ),
      .b_chan_t           (b_chan_t           ),
      .ar_chan_t          (ar_chan_t          ),
      .mst_r_chan_t       (mst_r_chan_t       ),
      .slv_r_chan_t       (slv_r_chan_t       ),
      .mst_port_axi_req_t (mst_port_axi_req_t ),
      .mst_port_axi_rsp_t (mst_port_axi_rsp_t ),
      .slv_port_axi_req_t (slv_port_axi_req_t ),
      .slv_port_axi_rsp_t (slv_port_axi_rsp_t )
    ) i_axi_dw_downsizer (
      .clk_i     (clk_i    ),
      .rst_ni    (rst_ni   ),
      // Slave interface
      .slv_req_i (slv_req_i),
      .slv_rsp_o (slv_rsp_o),
      // Master interface
      .mst_req_o (mst_req_o),
      .mst_rsp_i (mst_rsp_i)
    );
  end : gen_dw_downsize

endmodule : axi_dw_converter

// Interface wrapper

`include "axi/assign.svh"
`include "axi/typedef.svh"

module axi_dw_converter_intf #(
    parameter int unsigned AXI_ID_WIDTH            = 1,
    parameter int unsigned AXI_ADDR_WIDTH          = 1,
    parameter int unsigned AXI_SLV_PORT_DATA_WIDTH = 8,
    parameter int unsigned AXI_MST_PORT_DATA_WIDTH = 8,
    parameter int unsigned AXI_USER_WIDTH          = 0,
    parameter int unsigned AXI_MAX_READS           = 8
  ) (
    input          logic clk_i,
    input          logic rst_ni,
    AXI_BUS.Slave        slv,
    AXI_BUS.Master       mst
  );

  typedef logic [AXI_ID_WIDTH-1:0] id_t                   ;
  typedef logic [AXI_ADDR_WIDTH-1:0] addr_t               ;
  typedef logic [AXI_MST_PORT_DATA_WIDTH-1:0] mst_data_t  ;
  typedef logic [AXI_MST_PORT_DATA_WIDTH/8-1:0] mst_strb_t;
  typedef logic [AXI_SLV_PORT_DATA_WIDTH-1:0] slv_data_t  ;
  typedef logic [AXI_SLV_PORT_DATA_WIDTH/8-1:0] slv_strb_t;
  typedef logic [AXI_USER_WIDTH-1:0] user_t               ;
  `AXI_TYPEDEF_AW_CHAN_T(aw_chan_t, addr_t, id_t, user_t)
  `AXI_TYPEDEF_W_CHAN_T(mst_w_chan_t, mst_data_t, mst_strb_t, user_t)
  `AXI_TYPEDEF_W_CHAN_T(slv_w_chan_t, slv_data_t, slv_strb_t, user_t)
  `AXI_TYPEDEF_B_CHAN_T(b_chan_t, id_t, user_t)
  `AXI_TYPEDEF_AR_CHAN_T(ar_chan_t, addr_t, id_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(mst_r_chan_t, mst_data_t, id_t, user_t)
  `AXI_TYPEDEF_R_CHAN_T(slv_r_chan_t, slv_data_t, id_t, user_t)
  `AXI_TYPEDEF_REQ_T(mst_port_axi_req_t, aw_chan_t, mst_w_chan_t, ar_chan_t)
  `AXI_TYPEDEF_RSP_T(mst_port_axi_rsp_t, b_chan_t, mst_r_chan_t)
  `AXI_TYPEDEF_REQ_T(slv_port_axi_req_t, aw_chan_t, slv_w_chan_t, ar_chan_t)
  `AXI_TYPEDEF_RSP_T(slv_port_axi_rsp_t, b_chan_t, slv_r_chan_t)

  slv_port_axi_req_t slv_req;
  slv_port_axi_rsp_t slv_rsp;
  mst_port_axi_req_t mst_req;
  mst_port_axi_rsp_t mst_rsp;

  `AXI_ASSIGN_TO_REQ(slv_req, slv)
  `AXI_ASSIGN_FROM_RSP(slv, slv_rsp)

  `AXI_ASSIGN_FROM_REQ(mst, mst_req)
  `AXI_ASSIGN_TO_RSP(mst_rsp, mst)

  axi_dw_converter #(
    .MaxReads           ( AXI_MAX_READS           ),
    .SlvPortDataWidth   ( AXI_SLV_PORT_DATA_WIDTH ),
    .MstPortDataWidth   ( AXI_MST_PORT_DATA_WIDTH ),
    .AddrWidth          ( AXI_ADDR_WIDTH          ),
    .IdWidth            ( AXI_ID_WIDTH            ),
    .aw_chan_t          ( aw_chan_t               ),
    .mst_w_chan_t       ( mst_w_chan_t            ),
    .slv_w_chan_t       ( slv_w_chan_t            ),
    .b_chan_t           ( b_chan_t                ),
    .ar_chan_t          ( ar_chan_t               ),
    .mst_r_chan_t       ( mst_r_chan_t            ),
    .slv_r_chan_t       ( slv_r_chan_t            ),
    .mst_port_axi_req_t ( mst_port_axi_req_t               ),
    .mst_port_axi_rsp_t ( mst_port_axi_rsp_t               ),
    .slv_port_axi_req_t ( slv_port_axi_req_t               ),
    .slv_port_axi_rsp_t ( slv_port_axi_rsp_t               )
  ) i_axi_dw_converter (
    .clk_i      ( clk_i    ),
    .rst_ni     ( rst_ni   ),
    // slave port
    .slv_req_i  ( slv_req  ),
    .slv_rsp_o ( slv_rsp ),
    // master port
    .mst_req_o  ( mst_req  ),
    .mst_rsp_i ( mst_rsp )
  );

endmodule : axi_dw_converter_intf
